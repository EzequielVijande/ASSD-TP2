BZh91AY&SY�r 3߀Py���g߰����P��'s� �OS �&F  h�h �����4 � F@�@ h�"j��&��!�!�i 9�&& &#4���d�#�&F�&�1I�f�z�M �i�� -��@2E��|��b`����m�B��=L(4aW&s�p��H6˰@�!k�M�D�(�U�=[�
 �
1ֶ�$(jd�2�P3P���%L��M>�6{�d��bc��w˭x��}�^`���9=�%3���G���HH�:A�t �{����v�/�"L���G-8�,H���-:���ײ�Z�s$�Hq5��R��0{ɟ*��L '�AJc��pn&-@H,�`�P0�/&�b�Q�����J�c�]����_$��K.�'��-)�*���2�Y�5�4�
au�`�0n.Α�>���-���@a�d��3�f�?�[�c4�����X>:���QG�sAa�U�H(��_�9�*SYb�ߛ��d����p�|Ip����	XEG.2(ǒ�;�
8�Sb�E�@�fxy!M�I�M�>�_ю�0�gD�"pu��C[J'� Yh����p[���խnߤ�n"��B�""���&�b͜�IH?Y�w ���m[(���,��#
@�	��f6��Ao��Q
�d�	c$>��a�Md*�5�N"���ȓ�P��[{�!��a �/�{.-��'��'��}�� �^m#7i�ap��\��� ;�p3���Z)3�{h���H���79t�r1����l��	uӸ�7�T�[w�5��T�e}R;5�5�超B��h8Q#�g� Fa.�je!��f�c:�V~�����$]�ʮ?�w$S�		q0� 