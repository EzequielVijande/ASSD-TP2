BZh91AY&SYBu�� 5_�Py���g߰����P�� $�9�&& &#4���d�#hɉ�	���0 �`�0�"$�55?T<�Fi�='���  �4z�挘� ���F	� �D"`LJ���i������P2i�4hi���' 	���1� ����Ax��Cmi6�XB�lap�\®Y͔���i4I#����z)�`�6o�n׎N��|��j(�ԙXLn:bH4�:�R$�IJ.-
�f�!˗����;�a�PV�j�7YU��%��}�^���5�Dq�$niK�S�I^��{i]F�US�d�f�����;p�||~K�F4�塌i��m��<�Ύ�����)4�24��W'eo�s&����{J��P ���Y��3,�c��TM��ZٲlȬr���#����s4dAF�S��d����++`���gT�l���e��˱)+9�������U����Y� `*7�}Hx=A�1s�b�a���y
��ݨ�>���q�&b���D����^�C�����;o�/��� ��G�����o
1�� �y�s{�,H.��;ձ��I��Y�!IQ����I�KMM� ��/�����.DJ�9����W�D�>)�*H4��.r���b����t�E�0�)K�`��m�pL���u �[l�d4/�e&� �8OB+��p�[B%�418�@�.B�'OrT�C,��C�E�@�Q�R��*�y�	��;�}q�$=;9��'��i�0�y�0��ce�J�E�7�o+�
8� m9��N\0j�J!p��Z�RȀaŖs��lƓi},����h��)k;	ɣY
j�y�x��V�ݤ1/��D�2&�H���O��h�f�ւ��|�j12�&�)؎�{�|�t��.X�w$S�	'Xm`