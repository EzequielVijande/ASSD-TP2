BZh91AY&SY�U +_�Py���߰����P�t�ʀ�* j6��4i�Ƃz��z�2hɉ�	���0 �`�0�)��M��=M�ڞ���  4 �2b`b0#L1&L0H�@��T�d�4mL�������$(@ ��$	�_/�K�h(6�6�h�@�*�[
Uɝ��	���*�A�Z���͘	)F<��1��AV��ڐ�%�(��Z�!	)��,5����%`Z�����s��̓���\��:#pwv�� �&hN���$֝V:�v���/�6��J�Pω��������!	�D�I{�n��K0�!ȸD�2�9�_:̜�"����X�u	��s���IE)֚�mOV)P��e
'�_ǲ���v�C�N�;Ѻα�>��ȹV���5�a;�n�}�ǈd\e�u������,W�002D���2��&��H�Tw��"�����bp�{O:�=�F����Y�E���OaA��6�*�c�0�Vi�H�����$���-�H�?d����ҳ�悎4ڴ��l��PS,�M�.Ê_#F�0Ј\H��?�ze��q�;�������!�^��Ս���K��3^J��
��V��z̀ŎF4��C�`���n�4��h����Fj@�	��3[L��a9��\��,d���BV�M�C�h"���Q��,M|,�����Ựb��%��F�^{�=C��߀l�w���RA�>�v����M�u����@O�����)��2; !��āUR%�%���0��M9�tL8�g�ǧ!UIE�d`_�6k3=َmz1f�&P(�,�/Ί�B �%ˢ�b��j5��c:�V~�����H�q�\��H�
�
��