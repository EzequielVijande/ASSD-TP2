BZh91AY&SY���J *߀Py���g߰����P�t��(V�%M#F��j��d@�����@�sFLL LFi�#ɀF	M
L� с� @ 4�101��&$HF��C$x�I��#h#	�#�cD�`� �`?ᄁ3������~��mi6�\!\�V
0��8m0Xt$#�+ǹ,X�i�!	S��p���H+u�ό*5���X�:ł.�IJ���Q�ǟ厙X.Lu���Ի��X�T�H����|��Ș�Bhq��QE�3�8I�4��i�f�B��8[����>������˅$�C��1�����>$:_*ED��STP'
Ļ�"�`�5y$0TkӘz�f���}�ȕ��Zگ��V;Be�׾���tD+��%F�Q�SH�DS�:�md�Z��oI���"ʯ�����,4CJ�WS kX���B �Pq��De���4��}C��*0�����,������ D���4�F�-8�*S���n\ �gJ��ߘDn"]]"R�� �5tTp��tʅ�ݽe<)#AMkHt��@b��C�������	u����i���@�����ͫYD�`ȸ X�����xAS� ��ʬ
�ޘZԚ�BA�g+�9��-&T��C�ΰ�ٺ�r��[��B�`���H4��h���d'��H��*}(�,ơ��h#�V�&M1�I��%n�!�!�u� �zZ1>�	��6S%�����]8��,��Y��>�Iٰ�H��o��^���{�\J�-3#�BX������Se����b�u�Zh��H�6&�3	 Ȗ٫('��rX�p�P@{fP(�ɤc�+�:KnU3��~����F04)Ֆ�������$_�gW��w$S�	�]Ġ